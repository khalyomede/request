module request

pub struct ValidationRule {
	pub:
		rule Rule [required]
		parameters string
}
