module request

pub enum Rule {
	required
	filled
	boolean
}
